module Processing_element_tb2();
    parameter N=3,N_WIDTH=2,IFMAP_SIZE_WIDTH=4,GLOBAL_BUFFER_ADDR_WIDTH=10,GLOBAL_BUFFER_DEPTH=1000,STRIDE_WIDTH=2,FILTER_SIZE_WIDTH=4,IFMAP_ADDR_WIDTH=5,IFMAP_DEPTH=60,
    FILTER_ADDR_WIDTH=4,FILTER_DEPTH=10,DATA_WIDTH=16,IFMAP_BUF_DEPTH=60,PSUM_BUF_DEPTH=60,FILTER_BUF_DEPTH=60,PSUM_ADDR_WIDTH=5,PSUM_DEPTH=60;
    reg clk=0,rst=1,Start=0;
    reg [1:0] mode=2;
    reg [STRIDE_WIDTH-1:0] stride=1;
    reg [FILTER_SIZE_WIDTH-1:0] filter_size=5;
    reg [IFMAP_SIZE_WIDTH-1:0] ifmap_size=10;
    wire Done;

    PE_generator#(.N(N),.N_WIDTH(N_WIDTH),.GLOBAL_BUFFER_ADDR_WIDTH(GLOBAL_BUFFER_ADDR_WIDTH),.GLOBAL_BUFFER_DEPTH(GLOBAL_BUFFER_DEPTH),.STRIDE_WIDTH(STRIDE_WIDTH),.IFMAP_SIZE_WIDTH(IFMAP_SIZE_WIDTH),
    .FILTER_SIZE_WIDTH(FILTER_SIZE_WIDTH),.IFMAP_ADDR_WIDTH(IFMAP_ADDR_WIDTH),.IFMAP_DEPTH(IFMAP_DEPTH),.PSUM_ADDR_WIDTH(PSUM_ADDR_WIDTH),.PSUM_DEPTH(PSUM_DEPTH),
    .FILTER_ADDR_WIDTH(FILTER_ADDR_WIDTH),.FILTER_DEPTH(FILTER_DEPTH),.DATA_WIDTH(DATA_WIDTH),.PSUM_BUF_DEPTH(PSUM_BUF_DEPTH),.FILTER_BUF_DEPTH(FILTER_BUF_DEPTH),
    .IFMAP_BUF_DEPTH(IFMAP_BUF_DEPTH))PE_gen(.clk(clk),.rst(rst),.Start(Start),.mode(mode),.Done(Done),.stride(stride),.filter_size(filter_size),.ifmap_size(ifmap_size));

    always begin #19;clk=~clk;end
    initial begin
        #38;
        #38; rst=1'b0;
        #38; Start = 1'b1;
        #38; Start = 1'b0;
        #38000;
        $stop;
    end
endmodule